module mygate(input [0:0] a, input [0:0] b, output [0:0] c);

    assign c = a&b;

endmodule